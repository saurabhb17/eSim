* /home/ash98/eSim-Workspace/74LS32-test/74LS32-test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed Jan 15 20:34:15 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  in1 GND pulse		
v2  in2 GND pulse		
R1  in1 Net-_R1-Pad2_ 1k		
R3  in2 Net-_R3-Pad2_ 1k		
U1  in1 plot_v1		
U2  in2 plot_v1		
R2  out GND 1k		
U3  out plot_v1		
X1  Net-_R1-Pad2_ Net-_R3-Pad2_ out ? ? ? GND ? ? ? ? ? ? Net-_X1-Pad14_ eSim_74LS32		
v3  Net-_X1-Pad14_ GND DC		

.end
