* /home/ash98/eSim-Workspace/74LS00-test/74LS00-test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Jan 14 15:26:34 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  In1 Net-_R1-Pad2_ 1k		
R2  In2 Net-_R2-Pad2_ 1k		
v1  In1 GND pulse		
v2  In2 GND pulse		
U1  In1 plot_v1		
U2  In2 plot_v1		
v3  Net-_X1-Pad14_ GND DC		
R3  out GND 1k		
U3  out plot_v1		
X1  Net-_R1-Pad2_ Net-_R2-Pad2_ out ? ? ? GND ? ? ? ? ? ? Net-_X1-Pad14_ eSim_74LS00		

.end
