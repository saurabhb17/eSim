* /home/ash98/eSim-Workspace/74LS86-test/74LS86-test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu Jan 16 11:18:09 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  in1 in2 out ? ? ? GND ? ? ? ? ? ? Net-_X1-Pad14_ eSim_74LS86		
v1  in1 GND pulse		
v2  in2 GND pulse		
R1  out GND 1k		
v3  Net-_X1-Pad14_ GND DC		
U1  in1 plot_v1		
U2  in2 plot_v1		
U3  out plot_v1		

.end
