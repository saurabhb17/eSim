* /home/saurabh/Desktop/eSim/Examples/RC/RC.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat Feb  8 15:27:52 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
C1  out GND 1u		
R1  in out 1k		
U1  out plot_log		
U2  out plot_phase		
v1  in GND AC		

.end
