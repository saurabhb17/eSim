* /home/saurabh/Desktop/eSim/src/SubcircuitLibrary/74ls04/74ls04.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Jan 28 11:48:53 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_D1-Pad2_ Net-_D1-Pad1_ Net-_R1-Pad1_ Net-_Q4-Pad1_ PORT		
D2  Net-_D2-Pad1_ Net-_D1-Pad2_ eSim_Schottky		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Schottky		
Q1  Net-_D3-Pad2_ Net-_D2-Pad1_ Net-_Q1-Pad3_ eSim_NPN		
R2  Net-_D2-Pad1_ Net-_Q1-Pad3_ 12k		
R3  Net-_Q1-Pad3_ Net-_Q2-Pad2_ 1.5k		
Q2  Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_D1-Pad1_ eSim_NPN		
R5  Net-_Q1-Pad3_ Net-_Q2-Pad1_ 3k		
Q4  Net-_Q4-Pad1_ Net-_Q1-Pad3_ Net-_D1-Pad1_ eSim_NPN		
R1  Net-_R1-Pad1_ Net-_D2-Pad1_ 20k		
R4  Net-_R1-Pad1_ Net-_D3-Pad2_ 8k		
Q3  Net-_Q3-Pad1_ Net-_D3-Pad2_ Net-_D3-Pad1_ eSim_NPN		
R6  Net-_R1-Pad1_ Net-_Q3-Pad1_ 120		
D3  Net-_D3-Pad1_ Net-_D3-Pad2_ eSim_Schottky		
Q5  Net-_Q3-Pad1_ Net-_D3-Pad1_ Net-_Q4-Pad1_ eSim_NPN		
D4  Net-_D4-Pad1_ Net-_D3-Pad2_ eSim_Schottky		
R7  Net-_D3-Pad1_ Net-_D4-Pad1_ 4k		

.end
