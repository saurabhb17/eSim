* /home/ash98/Downloads/eSim-1.1.3/src/SubcircuitLibrary/3_and/3_and.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed Jan 15 16:55:49 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U2-Pad3_ d_and		
U3  Net-_U2-Pad3_ Net-_U3-Pad2_ Net-_U1-Pad4_ d_and		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ PORT		
U4  Net-_U1-Pad3_ Net-_U1-Pad3_ Net-_U3-Pad2_ d_and		

.end
